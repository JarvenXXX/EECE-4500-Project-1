*inverter

*declare parameters
.param plen = 70n
.param nlen = 70n
.param pwid = 220n
.param nwid = 130n
.param ptox = 1.95n
.param ntox = 1.85n

.subckt inverter in out plen=70n nlen=70n pwid=220n nwid=130n ptox=1.95n ntox=1.85n
M1 out in vdd vdd tp L=plen W=pwid
+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u
M2 out in vss vss tn L=nlen W=nwid
+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u

*BSIM 4.8.2 models
.model tp pmos level=54 version=4.8.2 toxp=ptox
.model tn nmos level=54 version=4.8.2 toxp=ntox

.ends inverter
